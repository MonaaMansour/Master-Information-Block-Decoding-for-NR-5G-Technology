module RateMatch (
    output reg [6 -1:0] mem_write_addr_r,
    output reg [2 -1:0] mem_llr_slct_r,
    output reg          llr_done_r,
    output reg          mem_1_w_enable_r,
    output reg          mem_2_w_enable_r,
    input wire          in_vld,
    input wire          clk,
    input wire          rst
);

reg [9:0] mem_write_addr;
reg [9:0] lut_read_addr_r;
reg [9:0] lut_read_addr;
reg       llr_done;
wire      mem_1_w_enable;
wire      mem_2_w_enable;


always @(posedge clk or negedge rst) begin
    if (!rst) begin
        mem_write_addr_r <= 'd0;
        lut_read_addr_r  <= 'd0;
        llr_done_r       <= 'd0;
        mem_1_w_enable_r <= 'd0;
        mem_2_w_enable_r <= 'd0;
        mem_llr_slct_r   <= 'd0;
    end
    else begin
        mem_write_addr_r <= mem_write_addr[7:2];
        mem_llr_slct_r   <= mem_write_addr[1:0];
        llr_done_r       <= llr_done;
        mem_1_w_enable_r <= mem_1_w_enable; 
        mem_2_w_enable_r <= mem_2_w_enable; 
        if(in_vld) begin
            lut_read_addr_r <= lut_read_addr;
        end
        
    end
end

assign  mem_1_w_enable  = in_vld && !mem_write_addr[8] && !mem_write_addr[9]; //mem_write_addr[8] to select between 2 rams
assign  mem_2_w_enable  = in_vld &&  mem_write_addr[8] && !mem_write_addr[9]; //mem_write_addr[9] to decide whether the input will be stored or ignored

always @(*) begin
    llr_done = 1'b0;
    lut_read_addr = lut_read_addr_r + 'd1;


    if (lut_read_addr_r == 'd863) begin
        llr_done = 1'b1;
        lut_read_addr = 'd0;
    end

    ///////////////LUT////////////////
    case (lut_read_addr_r)
        'd0   : mem_write_addr = 'd0;
        'd1   : mem_write_addr = 'd42;
        'd2   : mem_write_addr = 'd83;
        'd3   : mem_write_addr = 'd123;
        'd4   : mem_write_addr = 'd146;
        'd5   : mem_write_addr = 'd168;
        'd6   : mem_write_addr = 'd189;
        'd7   : mem_write_addr = 'd321;
        'd8   : mem_write_addr = 'd340;
        'd9   : mem_write_addr = 'd358;
        'd10  : mem_write_addr = 'd375;
        'd11  : mem_write_addr = 'd407;
        'd12  : mem_write_addr = 'd454;
        'd13  : mem_write_addr = 'd468;
        'd14  : mem_write_addr = 'd497;
        'd15  : mem_write_addr = 'd512;
        'd16  : mem_write_addr = 'd512;
        'd17  : mem_write_addr = 'd512;
        'd18  : mem_write_addr = 'd512;
        'd19  : mem_write_addr = 'd512;
        'd20  : mem_write_addr = 'd512;
        'd21  : mem_write_addr = 'd512;
        'd22  : mem_write_addr = 'd512;
        'd23  : mem_write_addr = 'd512;
        'd24  : mem_write_addr = 'd512;
        'd25  : mem_write_addr = 'd512;
        'd26  : mem_write_addr = 'd512;
        'd27  : mem_write_addr = 'd512;
        'd28  : mem_write_addr = 'd512;
        'd29  : mem_write_addr = 'd512;
        'd30  : mem_write_addr = 'd512;
        'd31  : mem_write_addr = 'd512;
        'd32  : mem_write_addr = 'd512;
        'd33  : mem_write_addr = 'd512;
        'd34  : mem_write_addr = 'd1;
        'd35  : mem_write_addr = 'd43;
        'd36  : mem_write_addr = 'd84;
        'd37  : mem_write_addr = 'd124;
        'd38  : mem_write_addr = 'd147;
        'd39  : mem_write_addr = 'd169;
        'd40  : mem_write_addr = 'd190;
        'd41  : mem_write_addr = 'd322;
        'd42  : mem_write_addr = 'd341;
        'd43  : mem_write_addr = 'd359;
        'd44  : mem_write_addr = 'd376;
        'd45  : mem_write_addr = 'd408;
        'd46  : mem_write_addr = 'd455;
        'd47  : mem_write_addr = 'd469;
        'd48  : mem_write_addr = 'd498;
        'd49  : mem_write_addr = 'd512;
        'd50  : mem_write_addr = 'd512;
        'd51  : mem_write_addr = 'd512;
        'd52  : mem_write_addr = 'd512;
        'd53  : mem_write_addr = 'd512;
        'd54  : mem_write_addr = 'd512;
        'd55  : mem_write_addr = 'd512;
        'd56  : mem_write_addr = 'd512;
        'd57  : mem_write_addr = 'd512;
        'd58  : mem_write_addr = 'd512;
        'd59  : mem_write_addr = 'd512;
        'd60  : mem_write_addr = 'd512;
        'd61  : mem_write_addr = 'd512;
        'd62  : mem_write_addr = 'd512;
        'd63  : mem_write_addr = 'd512;
        'd64  : mem_write_addr = 'd512;
        'd65  : mem_write_addr = 'd512;
        'd66  : mem_write_addr = 'd512;
        'd67  : mem_write_addr = 'd512;
        'd68  : mem_write_addr = 'd2;
        'd69  : mem_write_addr = 'd44;
        'd70  : mem_write_addr = 'd85;
        'd71  : mem_write_addr = 'd125;
        'd72  : mem_write_addr = 'd148;
        'd73  : mem_write_addr = 'd170;
        'd74  : mem_write_addr = 'd191;
        'd75  : mem_write_addr = 'd323;
        'd76  : mem_write_addr = 'd342;
        'd77  : mem_write_addr = 'd360;
        'd78  : mem_write_addr = 'd377;
        'd79  : mem_write_addr = 'd409;
        'd80  : mem_write_addr = 'd456;
        'd81  : mem_write_addr = 'd470;
        'd82  : mem_write_addr = 'd499;
        'd83  : mem_write_addr = 'd512;
        'd84  : mem_write_addr = 'd512;
        'd85  : mem_write_addr = 'd512;
        'd86  : mem_write_addr = 'd512;
        'd87  : mem_write_addr = 'd512;
        'd88  : mem_write_addr = 'd512;
        'd89  : mem_write_addr = 'd512;
        'd90  : mem_write_addr = 'd512;
        'd91  : mem_write_addr = 'd512;
        'd92  : mem_write_addr = 'd512;
        'd93  : mem_write_addr = 'd512;
        'd94  : mem_write_addr = 'd512;
        'd95  : mem_write_addr = 'd512;
        'd96  : mem_write_addr = 'd512;
        'd97  : mem_write_addr = 'd512;
        'd98  : mem_write_addr = 'd512;
        'd99  : mem_write_addr = 'd512;
        'd100 : mem_write_addr = 'd512;
        'd101 : mem_write_addr = 'd512;
        'd102 : mem_write_addr = 'd3;
        'd103 : mem_write_addr = 'd45;
        'd104 : mem_write_addr = 'd86;
        'd105 : mem_write_addr = 'd126;
        'd106 : mem_write_addr = 'd149;
        'd107 : mem_write_addr = 'd171;
        'd108 : mem_write_addr = 'd304;
        'd109 : mem_write_addr = 'd324;
        'd110 : mem_write_addr = 'd343;
        'd111 : mem_write_addr = 'd361;
        'd112 : mem_write_addr = 'd378;
        'd113 : mem_write_addr = 'd410;
        'd114 : mem_write_addr = 'd457;
        'd115 : mem_write_addr = 'd471;
        'd116 : mem_write_addr = 'd500;
        'd117 : mem_write_addr = 'd512;
        'd118 : mem_write_addr = 'd512;
        'd119 : mem_write_addr = 'd512;
        'd120 : mem_write_addr = 'd512;
        'd121 : mem_write_addr = 'd512;
        'd122 : mem_write_addr = 'd512;
        'd123 : mem_write_addr = 'd512;
        'd124 : mem_write_addr = 'd512;
        'd125 : mem_write_addr = 'd512;
        'd126 : mem_write_addr = 'd512;
        'd127 : mem_write_addr = 'd512;
        'd128 : mem_write_addr = 'd512;
        'd129 : mem_write_addr = 'd512;
        'd130 : mem_write_addr = 'd512;
        'd131 : mem_write_addr = 'd512;
        'd132 : mem_write_addr = 'd512;
        'd133 : mem_write_addr = 'd512;
        'd134 : mem_write_addr = 'd512;
        'd135 : mem_write_addr = 'd512;
        'd136 : mem_write_addr = 'd4;
        'd137 : mem_write_addr = 'd46;
        'd138 : mem_write_addr = 'd87;
        'd139 : mem_write_addr = 'd127;
        'd140 : mem_write_addr = 'd150;
        'd141 : mem_write_addr = 'd172;
        'd142 : mem_write_addr = 'd305;
        'd143 : mem_write_addr = 'd325;
        'd144 : mem_write_addr = 'd344;
        'd145 : mem_write_addr = 'd362;
        'd146 : mem_write_addr = 'd379;
        'd147 : mem_write_addr = 'd411;
        'd148 : mem_write_addr = 'd458;
        'd149 : mem_write_addr = 'd472;
        'd150 : mem_write_addr = 'd501;
        'd151 : mem_write_addr = 'd512;
        'd152 : mem_write_addr = 'd512;
        'd153 : mem_write_addr = 'd512;
        'd154 : mem_write_addr = 'd512;
        'd155 : mem_write_addr = 'd512;
        'd156 : mem_write_addr = 'd512;
        'd157 : mem_write_addr = 'd512;
        'd158 : mem_write_addr = 'd512;
        'd159 : mem_write_addr = 'd512;
        'd160 : mem_write_addr = 'd512;
        'd161 : mem_write_addr = 'd512;
        'd162 : mem_write_addr = 'd512;
        'd163 : mem_write_addr = 'd512;
        'd164 : mem_write_addr = 'd512;
        'd165 : mem_write_addr = 'd512;
        'd166 : mem_write_addr = 'd512;
        'd167 : mem_write_addr = 'd512;
        'd168 : mem_write_addr = 'd512;
        'd169 : mem_write_addr = 'd512;//
        'd170 : mem_write_addr = 'd5;
        'd171 : mem_write_addr = 'd47;
        'd172 : mem_write_addr = 'd88;
        'd173 : mem_write_addr = 'd128;
        'd174 : mem_write_addr = 'd151;
        'd175 : mem_write_addr = 'd173;
        'd176 : mem_write_addr = 'd306;
        'd177 : mem_write_addr = 'd326;
        'd178 : mem_write_addr = 'd345;
        'd179 : mem_write_addr = 'd363;//
        'd180 : mem_write_addr = 'd380;
        'd181 : mem_write_addr = 'd412;
        'd182 : mem_write_addr = 'd459;
        'd183 : mem_write_addr = 'd473;
        'd184 : mem_write_addr = 'd502;
        'd185 : mem_write_addr = 'd512;
        'd186 : mem_write_addr = 'd512;
        'd187 : mem_write_addr = 'd512;
        'd188 : mem_write_addr = 'd512;
        'd189 : mem_write_addr = 'd512;//
        'd190 : mem_write_addr = 'd512;
        'd191 : mem_write_addr = 'd512;
        'd192 : mem_write_addr = 'd512;
        'd193 : mem_write_addr = 'd512;
        'd194 : mem_write_addr = 'd512;
        'd195 : mem_write_addr = 'd512;
        'd196 : mem_write_addr = 'd512;
        'd197 : mem_write_addr = 'd512;
        'd198 : mem_write_addr = 'd512;
        'd199 : mem_write_addr = 'd512;//
        'd200 : mem_write_addr = 'd512;
        'd201 : mem_write_addr = 'd512;
        'd202 : mem_write_addr = 'd512;
        'd203 : mem_write_addr = 'd512;
        'd204 : mem_write_addr = 'd6;
        'd205 : mem_write_addr = 'd64;
        'd206 : mem_write_addr = 'd89;
        'd207 : mem_write_addr = 'd129;
        'd208 : mem_write_addr = 'd152;
        'd209 : mem_write_addr = 'd174;//
        'd210 : mem_write_addr = 'd307;
        'd211 : mem_write_addr = 'd327;
        'd212 : mem_write_addr = 'd346;
        'd213 : mem_write_addr = 'd364;
        'd214 : mem_write_addr = 'd381;
        'd215 : mem_write_addr = 'd413;
        'd216 : mem_write_addr = 'd460;
        'd217 : mem_write_addr = 'd474;
        'd218 : mem_write_addr = 'd503;
        'd219 : mem_write_addr = 'd512;//
        'd220 : mem_write_addr = 'd512;
        'd221 : mem_write_addr = 'd512;
        'd222 : mem_write_addr = 'd512;
        'd223 : mem_write_addr = 'd512;
        'd224 : mem_write_addr = 'd512;
        'd225 : mem_write_addr = 'd512;
        'd226 : mem_write_addr = 'd512;
        'd227 : mem_write_addr = 'd512;
        'd228 : mem_write_addr = 'd512;
        'd229 : mem_write_addr = 'd512;//
        'd230 : mem_write_addr = 'd512;
        'd231 : mem_write_addr = 'd512;
        'd232 : mem_write_addr = 'd512;
        'd233 : mem_write_addr = 'd512;
        'd234 : mem_write_addr = 'd512;
        'd235 : mem_write_addr = 'd512;
        'd236 : mem_write_addr = 'd512;
        'd237 : mem_write_addr = 'd7;
        'd238 : mem_write_addr = 'd65;
        'd239 : mem_write_addr = 'd90;//
        'd240 : mem_write_addr = 'd130;
        'd241 : mem_write_addr = 'd153;
        'd242 : mem_write_addr = 'd175;
        'd243 : mem_write_addr = 'd308;
        'd244 : mem_write_addr = 'd328;
        'd245 : mem_write_addr = 'd347;
        'd246 : mem_write_addr = 'd365;
        'd247 : mem_write_addr = 'd382;
        'd248 : mem_write_addr = 'd414;
        'd249 : mem_write_addr = 'd461;//
        'd250 : mem_write_addr = 'd475;
        'd251 : mem_write_addr = 'd504;
        'd252 : mem_write_addr = 'd512;
        'd253 : mem_write_addr = 'd512;
        'd254 : mem_write_addr = 'd512;
        'd255 : mem_write_addr = 'd512;
        'd256 : mem_write_addr = 'd512;
        'd257 : mem_write_addr = 'd512;
        'd258 : mem_write_addr = 'd512;
        'd259 : mem_write_addr = 'd512;//
        'd260 : mem_write_addr = 'd512;
        'd261 : mem_write_addr = 'd512;
        'd262 : mem_write_addr = 'd512;
        'd263 : mem_write_addr = 'd512;
        'd264 : mem_write_addr = 'd512;
        'd265 : mem_write_addr = 'd512;
        'd266 : mem_write_addr = 'd512;
        'd267 : mem_write_addr = 'd512;
        'd268 : mem_write_addr = 'd512;
        'd269 : mem_write_addr = 'd512;//
        'd270 : mem_write_addr = 'd8;
        'd271 : mem_write_addr = 'd66;
        'd272 : mem_write_addr = 'd91;
        'd273 : mem_write_addr = 'd131;
        'd274 : mem_write_addr = 'd154;
        'd275 : mem_write_addr = 'd288;
        'd276 : mem_write_addr = 'd309;
        'd277 : mem_write_addr = 'd329;
        'd278 : mem_write_addr = 'd348;
        'd279 : mem_write_addr = 'd366;//
        'd280 : mem_write_addr = 'd383;
        'd281 : mem_write_addr = 'd415;
        'd282 : mem_write_addr = 'd462;
        'd283 : mem_write_addr = 'd476;
        'd284 : mem_write_addr = 'd505;
        'd285 : mem_write_addr = 'd512;
        'd286 : mem_write_addr = 'd512;
        'd287 : mem_write_addr = 'd512;
        'd288 : mem_write_addr = 'd512;
        'd289 : mem_write_addr = 'd512;//
        'd290 : mem_write_addr = 'd512;
        'd291 : mem_write_addr = 'd512;
        'd292 : mem_write_addr = 'd512;
        'd293 : mem_write_addr = 'd512;
        'd294 : mem_write_addr = 'd512;
        'd295 : mem_write_addr = 'd512;
        'd296 : mem_write_addr = 'd512;
        'd297 : mem_write_addr = 'd512;
        'd298 : mem_write_addr = 'd512;
        'd299 : mem_write_addr = 'd512;//
        'd300 : mem_write_addr = 'd512;
        'd301 : mem_write_addr = 'd512;
        'd302 : mem_write_addr = 'd512;
        'd303 : mem_write_addr = 'd9;
        'd304 : mem_write_addr = 'd67;
        'd305 : mem_write_addr = 'd92;
        'd306 : mem_write_addr = 'd132;
        'd307 : mem_write_addr = 'd155;
        'd308 : mem_write_addr = 'd289;
        'd309 : mem_write_addr = 'd310;//
        'd310 : mem_write_addr = 'd330;
        'd311 : mem_write_addr = 'd349;
        'd312 : mem_write_addr = 'd367;
        'd313 : mem_write_addr = 'd384;
        'd314 : mem_write_addr = 'd416;
        'd315 : mem_write_addr = 'd463;
        'd316 : mem_write_addr = 'd477;
        'd317 : mem_write_addr = 'd506;
        'd318 : mem_write_addr = 'd512;
        'd319 : mem_write_addr = 'd512;//
        'd320 : mem_write_addr = 'd512;
        'd321 : mem_write_addr = 'd512;
        'd322 : mem_write_addr = 'd512;
        'd323 : mem_write_addr = 'd512;
        'd324 : mem_write_addr = 'd512;
        'd325 : mem_write_addr = 'd512;
        'd326 : mem_write_addr = 'd512;
        'd327 : mem_write_addr = 'd512;
        'd328 : mem_write_addr = 'd512;
        'd329 : mem_write_addr = 'd512;//
        'd330 : mem_write_addr = 'd512;
        'd331 : mem_write_addr = 'd512;
        'd332 : mem_write_addr = 'd512;
        'd333 : mem_write_addr = 'd512;
        'd334 : mem_write_addr = 'd512;
        'd335 : mem_write_addr = 'd512;
        'd336 : mem_write_addr = 'd10;
        'd337 : mem_write_addr = 'd68;
        'd338 : mem_write_addr = 'd93;
        'd339 : mem_write_addr = 'd133;//
        'd340 : mem_write_addr = 'd156;
        'd341 : mem_write_addr = 'd290;
        'd342 : mem_write_addr = 'd311;
        'd343 : mem_write_addr = 'd331;
        'd344 : mem_write_addr = 'd350;
        'd345 : mem_write_addr = 'd240;
        'd346 : mem_write_addr = 'd385;
        'd347 : mem_write_addr = 'd417;
        'd348 : mem_write_addr = 'd432;
        'd349 : mem_write_addr = 'd478;//
        'd350 : mem_write_addr = 'd507;
        'd351 : mem_write_addr = 'd512;
        'd352 : mem_write_addr = 'd512;
        'd353 : mem_write_addr = 'd512;
        'd354 : mem_write_addr = 'd512;
        'd355 : mem_write_addr = 'd512;
        'd356 : mem_write_addr = 'd512;
        'd357 : mem_write_addr = 'd512;
        'd358 : mem_write_addr = 'd512;
        'd359 : mem_write_addr = 'd512;//
        'd360 : mem_write_addr = 'd512;
        'd361 : mem_write_addr = 'd512;
        'd362 : mem_write_addr = 'd512;
        'd363 : mem_write_addr = 'd512;
        'd364 : mem_write_addr = 'd512;
        'd365 : mem_write_addr = 'd512;
        'd366 : mem_write_addr = 'd512;
        'd367 : mem_write_addr = 'd512;
        'd368 : mem_write_addr = 'd11;
        'd369 : mem_write_addr = 'd69;//
        'd370 : mem_write_addr = 'd94;
        'd371 : mem_write_addr = 'd134;
        'd372 : mem_write_addr = 'd157;
        'd373 : mem_write_addr = 'd291;
        'd374 : mem_write_addr = 'd312;
        'd375 : mem_write_addr = 'd332;
        'd376 : mem_write_addr = 'd351;
        'd377 : mem_write_addr = 'd241;
        'd378 : mem_write_addr = 'd386;
        'd379 : mem_write_addr = 'd418;//
        'd380 : mem_write_addr = 'd433;
        'd381 : mem_write_addr = 'd479;
        'd382 : mem_write_addr = 'd508;
        'd383 : mem_write_addr = 'd512;
        'd384 : mem_write_addr = 'd512;
        'd385 : mem_write_addr = 'd512;
        'd386 : mem_write_addr = 'd512;
        'd387 : mem_write_addr = 'd512;
        'd388 : mem_write_addr = 'd512;
        'd389 : mem_write_addr = 'd512;//
        'd390 : mem_write_addr = 'd512;
        'd391 : mem_write_addr = 'd512;
        'd392 : mem_write_addr = 'd512;
        'd393 : mem_write_addr = 'd512;
        'd394 : mem_write_addr = 'd512;
        'd395 : mem_write_addr = 'd512;
        'd396 : mem_write_addr = 'd512;
        'd397 : mem_write_addr = 'd512;
        'd398 : mem_write_addr = 'd512;
        'd399 : mem_write_addr = 'd12;//
        'd400 : mem_write_addr = 'd70;
        'd401 : mem_write_addr = 'd95;
        'd402 : mem_write_addr = 'd135;
        'd403 : mem_write_addr = 'd158;
        'd404 : mem_write_addr = 'd292;
        'd405 : mem_write_addr = 'd313;
        'd406 : mem_write_addr = 'd333;
        'd407 : mem_write_addr = 'd224;
        'd408 : mem_write_addr = 'd242;
        'd409 : mem_write_addr = 'd387;//
        'd410 : mem_write_addr = 'd419;
        'd411 : mem_write_addr = 'd434;
        'd412 : mem_write_addr = 'd480;
        'd413 : mem_write_addr = 'd509;
        'd414 : mem_write_addr = 'd512;
        'd415 : mem_write_addr = 'd512;
        'd416 : mem_write_addr = 'd512;
        'd417 : mem_write_addr = 'd512;
        'd418 : mem_write_addr = 'd512;
        'd419 : mem_write_addr = 'd512;//
        'd420 : mem_write_addr = 'd512;
        'd421 : mem_write_addr = 'd512;
        'd422 : mem_write_addr = 'd512;
        'd423 : mem_write_addr = 'd512;
        'd424 : mem_write_addr = 'd512;
        'd425 : mem_write_addr = 'd512;
        'd426 : mem_write_addr = 'd512;
        'd427 : mem_write_addr = 'd512;
        'd428 : mem_write_addr = 'd512;
        'd429 : mem_write_addr = 'd13;//
        'd430 : mem_write_addr = 'd71;
        'd431 : mem_write_addr = 'd96;
        'd432 : mem_write_addr = 'd136;
        'd433 : mem_write_addr = 'd159;
        'd434 : mem_write_addr = 'd293;
        'd435 : mem_write_addr = 'd314;
        'd436 : mem_write_addr = 'd334;
        'd437 : mem_write_addr = 'd225;
        'd438 : mem_write_addr = 'd243;
        'd439 : mem_write_addr = 'd388;//
        'd440 : mem_write_addr = 'd420;
        'd441 : mem_write_addr = 'd435;
        'd442 : mem_write_addr = 'd481;
        'd443 : mem_write_addr = 'd510;
        'd444 : mem_write_addr = 'd512;
        'd445 : mem_write_addr = 'd512;
        'd446 : mem_write_addr = 'd512;
        'd447 : mem_write_addr = 'd512;
        'd448 : mem_write_addr = 'd512;
        'd449 : mem_write_addr = 'd512;//
        'd450 : mem_write_addr = 'd512;
        'd451 : mem_write_addr = 'd512;
        'd452 : mem_write_addr = 'd512;
        'd453 : mem_write_addr = 'd512;
        'd454 : mem_write_addr = 'd512;
        'd455 : mem_write_addr = 'd512;
        'd456 : mem_write_addr = 'd512;
        'd457 : mem_write_addr = 'd512;
        'd458 : mem_write_addr = 'd14;
        'd459 : mem_write_addr = 'd72;//
        'd460 : mem_write_addr = 'd97;
        'd461 : mem_write_addr = 'd137;
        'd462 : mem_write_addr = 'd272;
        'd463 : mem_write_addr = 'd294;
        'd464 : mem_write_addr = 'd315;
        'd465 : mem_write_addr = 'd335;
        'd466 : mem_write_addr = 'd226;
        'd467 : mem_write_addr = 'd244;
        'd468 : mem_write_addr = 'd389;
        'd469 : mem_write_addr = 'd421;//  
        'd470 : mem_write_addr = 'd436;
        'd471 : mem_write_addr = 'd482;
        'd472 : mem_write_addr = 'd511;
        'd473 : mem_write_addr = 'd512;
        'd474 : mem_write_addr = 'd512;
        'd475 : mem_write_addr = 'd512;
        'd476 : mem_write_addr = 'd512;
        'd477 : mem_write_addr = 'd512;
        'd478 : mem_write_addr = 'd512;
        'd479 : mem_write_addr = 'd512;//
        'd480 : mem_write_addr = 'd512;
        'd481 : mem_write_addr = 'd512;
        'd482 : mem_write_addr = 'd512;
        'd483 : mem_write_addr = 'd512;
        'd484 : mem_write_addr = 'd512;
        'd485 : mem_write_addr = 'd512;
        'd486 : mem_write_addr = 'd15;
        'd487 : mem_write_addr = 'd73;
        'd488 : mem_write_addr = 'd98;
        'd489 : mem_write_addr = 'd138;//
        'd490 : mem_write_addr = 'd273;
        'd491 : mem_write_addr = 'd295;
        'd492 : mem_write_addr = 'd316;
        'd493 : mem_write_addr = 'd208;
        'd494 : mem_write_addr = 'd227;
        'd495 : mem_write_addr = 'd245;
        'd496 : mem_write_addr = 'd390;
        'd497 : mem_write_addr = 'd422;
        'd498 : mem_write_addr = 'd437;
        'd499 : mem_write_addr = 'd483;//
        'd500 : mem_write_addr = 'd512;
        'd501 : mem_write_addr = 'd512;
        'd502 : mem_write_addr = 'd512;
        'd503 : mem_write_addr = 'd512;
        'd504 : mem_write_addr = 'd512;
        'd505 : mem_write_addr = 'd512;
        'd506 : mem_write_addr = 'd512;
        'd507 : mem_write_addr = 'd512;
        'd508 : mem_write_addr = 'd512;
        'd509 : mem_write_addr = 'd512;//
        'd510 : mem_write_addr = 'd512;
        'd511 : mem_write_addr = 'd512;
        'd512 : mem_write_addr = 'd512;
        'd513 : mem_write_addr = 'd16;
        'd514 : mem_write_addr = 'd74;
        'd515 : mem_write_addr = 'd99;
        'd516 : mem_write_addr = 'd139;
        'd517 : mem_write_addr = 'd274;
        'd518 : mem_write_addr = 'd296;
        'd519 : mem_write_addr = 'd317;//
        'd520 : mem_write_addr = 'd209;
        'd521 : mem_write_addr = 'd228;
        'd522 : mem_write_addr = 'd246;
        'd523 : mem_write_addr = 'd391;
        'd524 : mem_write_addr = 'd423;
        'd525 : mem_write_addr = 'd438;
        'd526 : mem_write_addr = 'd484;
        'd527 : mem_write_addr = 'd512;
        'd528 : mem_write_addr = 'd512;
        'd529 : mem_write_addr = 'd512;//
        'd530 : mem_write_addr = 'd512;
        'd531 : mem_write_addr = 'd512;
        'd532 : mem_write_addr = 'd512;
        'd533 : mem_write_addr = 'd512;
        'd534 : mem_write_addr = 'd512;
        'd535 : mem_write_addr = 'd512;
        'd536 : mem_write_addr = 'd512;
        'd537 : mem_write_addr = 'd512;
        'd538 : mem_write_addr = 'd512;
        'd539 : mem_write_addr = 'd17;//  
        'd540 : mem_write_addr = 'd75;
        'd541 : mem_write_addr = 'd100;
        'd542 : mem_write_addr = 'd140;
        'd543 : mem_write_addr = 'd275;
        'd544 : mem_write_addr = 'd297;
        'd545 : mem_write_addr = 'd318;
        'd546 : mem_write_addr = 'd210;
        'd547 : mem_write_addr = 'd229;
        'd548 : mem_write_addr = 'd247;
        'd549 : mem_write_addr = 'd392;//
        'd550 : mem_write_addr = 'd424;
        'd551 : mem_write_addr = 'd439;
        'd552 : mem_write_addr = 'd485;
        'd553 : mem_write_addr = 'd512;
        'd554 : mem_write_addr = 'd512;
        'd555 : mem_write_addr = 'd512;
        'd556 : mem_write_addr = 'd512;
        'd557 : mem_write_addr = 'd512;
        'd558 : mem_write_addr = 'd512;
        'd559 : mem_write_addr = 'd512;//
        'd560 : mem_write_addr = 'd512;
        'd561 : mem_write_addr = 'd512;
        'd562 : mem_write_addr = 'd512;
        'd563 : mem_write_addr = 'd512;
        'd564 : mem_write_addr = 'd18;
        'd565 : mem_write_addr = 'd76;
        'd566 : mem_write_addr = 'd101;
        'd567 : mem_write_addr = 'd141;
        'd568 : mem_write_addr = 'd276;
        'd569 : mem_write_addr = 'd298;//
        'd570 : mem_write_addr = 'd319;
        'd571 : mem_write_addr = 'd211;
        'd572 : mem_write_addr = 'd230;
        'd573 : mem_write_addr = 'd248;
        'd574 : mem_write_addr = 'd393;
        'd575 : mem_write_addr = 'd425;
        'd576 : mem_write_addr = 'd440;
        'd577 : mem_write_addr = 'd486;
        'd578 : mem_write_addr = 'd512;
        'd579 : mem_write_addr = 'd512;// 
        'd580 : mem_write_addr = 'd512;
        'd581 : mem_write_addr = 'd512;
        'd582 : mem_write_addr = 'd512;
        'd583 : mem_write_addr = 'd512;
        'd584 : mem_write_addr = 'd512;
        'd585 : mem_write_addr = 'd512;
        'd586 : mem_write_addr = 'd512;
        'd587 : mem_write_addr = 'd512;
        'd588 : mem_write_addr = 'd19;
        'd589 : mem_write_addr = 'd77;//
        'd590 : mem_write_addr = 'd102;
        'd591 : mem_write_addr = 'd142;
        'd592 : mem_write_addr = 'd277;
        'd593 : mem_write_addr = 'd299;
        'd594 : mem_write_addr = 'd192;
        'd595 : mem_write_addr = 'd212;
        'd596 : mem_write_addr = 'd231;
        'd597 : mem_write_addr = 'd249;
        'd598 : mem_write_addr = 'd394;
        'd599 : mem_write_addr = 'd426;//
        'd600 : mem_write_addr = 'd441;
        'd601 : mem_write_addr = 'd487;
        'd602 : mem_write_addr = 'd512;
        'd603 : mem_write_addr = 'd512;
        'd604 : mem_write_addr = 'd512;
        'd605 : mem_write_addr = 'd512;
        'd606 : mem_write_addr = 'd512;
        'd607 : mem_write_addr = 'd512;
        'd608 : mem_write_addr = 'd512;
        'd609 : mem_write_addr = 'd512;//
        'd610 : mem_write_addr = 'd512;
        'd611 : mem_write_addr = 'd20;
        'd612 : mem_write_addr = 'd78;
        'd613 : mem_write_addr = 'd103;
        'd614 : mem_write_addr = 'd143;
        'd615 : mem_write_addr = 'd278;
        'd616 : mem_write_addr = 'd300;
        'd617 : mem_write_addr = 'd193;
        'd618 : mem_write_addr = 'd213;
        'd619 : mem_write_addr = 'd232;// 
        'd620 : mem_write_addr = 'd250;
        'd621 : mem_write_addr = 'd395;
        'd622 : mem_write_addr = 'd427;
        'd623 : mem_write_addr = 'd442;
        'd624 : mem_write_addr = 'd488;
        'd625 : mem_write_addr = 'd512;
        'd626 : mem_write_addr = 'd512;
        'd627 : mem_write_addr = 'd512;
        'd628 : mem_write_addr = 'd512;
        'd629 : mem_write_addr = 'd512;//
        'd630 : mem_write_addr = 'd512;
        'd631 : mem_write_addr = 'd512;
        'd632 : mem_write_addr = 'd512;
        'd633 : mem_write_addr = 'd21;
        'd634 : mem_write_addr = 'd79;
        'd635 : mem_write_addr = 'd104;
        'd636 : mem_write_addr = 'd256;
        'd637 : mem_write_addr = 'd279;
        'd638 : mem_write_addr = 'd301;
        'd639 : mem_write_addr = 'd194;//
        'd640 : mem_write_addr = 'd214;
        'd641 : mem_write_addr = 'd233;
        'd642 : mem_write_addr = 'd251;
        'd643 : mem_write_addr = 'd396;
        'd644 : mem_write_addr = 'd428;
        'd645 : mem_write_addr = 'd443;
        'd646 : mem_write_addr = 'd489;
        'd647 : mem_write_addr = 'd512;
        'd648 : mem_write_addr = 'd512;
        'd649 : mem_write_addr = 'd512;//
        'd650 : mem_write_addr = 'd512;
        'd651 : mem_write_addr = 'd512;
        'd652 : mem_write_addr = 'd512;
        'd653 : mem_write_addr = 'd512;
        'd654 : mem_write_addr = 'd22;
        'd655 : mem_write_addr = 'd48;
        'd656 : mem_write_addr = 'd105;
        'd657 : mem_write_addr = 'd257;
        'd658 : mem_write_addr = 'd280;
        'd659 : mem_write_addr = 'd302;// 
        'd660 : mem_write_addr = 'd195;
        'd661 : mem_write_addr = 'd215;
        'd662 : mem_write_addr = 'd234;
        'd663 : mem_write_addr = 'd252;
        'd664 : mem_write_addr = 'd397;
        'd665 : mem_write_addr = 'd429;
        'd666 : mem_write_addr = 'd444;
        'd667 : mem_write_addr = 'd490;
        'd668 : mem_write_addr = 'd512;
        'd669 : mem_write_addr = 'd512;//
        'd670 : mem_write_addr = 'd512;
        'd671 : mem_write_addr = 'd512;
        'd672 : mem_write_addr = 'd512;
        'd673 : mem_write_addr = 'd512;
        'd674 : mem_write_addr = 'd23;
        'd675 : mem_write_addr = 'd49;
        'd676 : mem_write_addr = 'd106;
        'd677 : mem_write_addr = 'd258;
        'd678 : mem_write_addr = 'd281;
        'd679 : mem_write_addr = 'd303;// 
        'd680 : mem_write_addr = 'd196;
        'd681 : mem_write_addr = 'd216;
        'd682 : mem_write_addr = 'd235;
        'd683 : mem_write_addr = 'd253;
        'd684 : mem_write_addr = 'd398;
        'd685 : mem_write_addr = 'd430;
        'd686 : mem_write_addr = 'd445;
        'd687 : mem_write_addr = 'd491;
        'd688 : mem_write_addr = 'd512;
        'd689 : mem_write_addr = 'd512;//
        'd690 : mem_write_addr = 'd512;
        'd691 : mem_write_addr = 'd512;
        'd692 : mem_write_addr = 'd512;
        'd693 : mem_write_addr = 'd24;
        'd694 : mem_write_addr = 'd50;
        'd695 : mem_write_addr = 'd107;
        'd696 : mem_write_addr = 'd259;
        'd697 : mem_write_addr = 'd282;
        'd698 : mem_write_addr = 'd176;
        'd699 : mem_write_addr = 'd197;//
        'd700 : mem_write_addr = 'd217;
        'd701 : mem_write_addr = 'd236;
        'd702 : mem_write_addr = 'd254;
        'd703 : mem_write_addr = 'd399;
        'd704 : mem_write_addr = 'd431;
        'd705 : mem_write_addr = 'd446;
        'd706 : mem_write_addr = 'd492;
        'd707 : mem_write_addr = 'd512;
        'd708 : mem_write_addr = 'd512;
        'd709 : mem_write_addr = 'd512;//
        'd710 : mem_write_addr = 'd512;
        'd711 : mem_write_addr = 'd25;
        'd712 : mem_write_addr = 'd51;
        'd713 : mem_write_addr = 'd108;
        'd714 : mem_write_addr = 'd260;
        'd715 : mem_write_addr = 'd283;
        'd716 : mem_write_addr = 'd177;
        'd717 : mem_write_addr = 'd198;
        'd718 : mem_write_addr = 'd218;
        'd719 : mem_write_addr = 'd237;// 
        'd720 : mem_write_addr = 'd255;
        'd721 : mem_write_addr = 'd400;
        'd722 : mem_write_addr = 'd448;
        'd723 : mem_write_addr = 'd447;
        'd724 : mem_write_addr = 'd493;
        'd725 : mem_write_addr = 'd512;
        'd726 : mem_write_addr = 'd512;
        'd727 : mem_write_addr = 'd512;
        'd728 : mem_write_addr = 'd26;
        'd729 : mem_write_addr = 'd52;//
        'd730 : mem_write_addr = 'd109;
        'd731 : mem_write_addr = 'd261;
        'd732 : mem_write_addr = 'd284;
        'd733 : mem_write_addr = 'd178;
        'd734 : mem_write_addr = 'd199;
        'd735 : mem_write_addr = 'd219;
        'd736 : mem_write_addr = 'd238;
        'd737 : mem_write_addr = 'd368;
        'd738 : mem_write_addr = 'd401;
        'd739 : mem_write_addr = 'd449;// 
        'd740 : mem_write_addr = 'd464;
        'd741 : mem_write_addr = 'd494;
        'd742 : mem_write_addr = 'd512;
        'd743 : mem_write_addr = 'd512;
        'd744 : mem_write_addr = 'd27;
        'd745 : mem_write_addr = 'd53;
        'd746 : mem_write_addr = 'd110;
        'd747 : mem_write_addr = 'd262;
        'd748 : mem_write_addr = 'd285;
        'd749 : mem_write_addr = 'd179;//
        'd750 : mem_write_addr = 'd200;
        'd751 : mem_write_addr = 'd220;
        'd752 : mem_write_addr = 'd239;
        'd753 : mem_write_addr = 'd369;
        'd754 : mem_write_addr = 'd402;
        'd755 : mem_write_addr = 'd450;
        'd756 : mem_write_addr = 'd465;
        'd757 : mem_write_addr = 'd495;
        'd758 : mem_write_addr = 'd512;
        'd759 : mem_write_addr = 'd28;//
        'd760 : mem_write_addr = 'd54;
        'd761 : mem_write_addr = 'd111;
        'd762 : mem_write_addr = 'd263;
        'd763 : mem_write_addr = 'd286;
        'd764 : mem_write_addr = 'd180;
        'd765 : mem_write_addr = 'd201;
        'd766 : mem_write_addr = 'd221;
        'd767 : mem_write_addr = 'd352;
        'd768 : mem_write_addr = 'd370;
        'd769 : mem_write_addr = 'd403;//
        'd770 : mem_write_addr = 'd451;
        'd771 : mem_write_addr = 'd466;
        'd772 : mem_write_addr = 'd496;
        'd773 : mem_write_addr = 'd29;
        'd774 : mem_write_addr = 'd55;
        'd775 : mem_write_addr = 'd112;
        'd776 : mem_write_addr = 'd264;
        'd777 : mem_write_addr = 'd287;
        'd778 : mem_write_addr = 'd181;
        'd779 : mem_write_addr = 'd202;// 
        'd780 : mem_write_addr = 'd222;
        'd781 : mem_write_addr = 'd353;
        'd782 : mem_write_addr = 'd371;
        'd783 : mem_write_addr = 'd404;
        'd784 : mem_write_addr = 'd452;
        'd785 : mem_write_addr = 'd467;
        'd786 : mem_write_addr = 'd30;
        'd787 : mem_write_addr = 'd56;
        'd788 : mem_write_addr = 'd113;
        'd789 : mem_write_addr = 'd265;//
        'd790 : mem_write_addr = 'd160;
        'd791 : mem_write_addr = 'd182;
        'd792 : mem_write_addr = 'd203;
        'd793 : mem_write_addr = 'd223;
        'd794 : mem_write_addr = 'd354;
        'd795 : mem_write_addr = 'd372;
        'd796 : mem_write_addr = 'd405;
        'd797 : mem_write_addr = 'd453;
        'd798 : mem_write_addr = 'd31;
        'd799 : mem_write_addr = 'd57;// 
        'd800 : mem_write_addr = 'd114;
        'd801 : mem_write_addr = 'd266;
        'd802 : mem_write_addr = 'd161;
        'd803 : mem_write_addr = 'd183;
        'd804 : mem_write_addr = 'd204;
        'd805 : mem_write_addr = 'd336;
        'd806 : mem_write_addr = 'd355;
        'd807 : mem_write_addr = 'd373;
        'd808 : mem_write_addr = 'd406;
        'd809 : mem_write_addr = 'd32;//
        'd810 : mem_write_addr = 'd58;
        'd811 : mem_write_addr = 'd115;
        'd812 : mem_write_addr = 'd267;
        'd813 : mem_write_addr = 'd162;
        'd814 : mem_write_addr = 'd184;
        'd815 : mem_write_addr = 'd205;
        'd816 : mem_write_addr = 'd337;
        'd817 : mem_write_addr = 'd356;
        'd818 : mem_write_addr = 'd374;
        'd819 : mem_write_addr = 'd33;//
        'd820 : mem_write_addr = 'd59;
        'd821 : mem_write_addr = 'd116;
        'd822 : mem_write_addr = 'd268;
        'd823 : mem_write_addr = 'd163;
        'd824 : mem_write_addr = 'd185;
        'd825 : mem_write_addr = 'd206;
        'd826 : mem_write_addr = 'd338;
        'd827 : mem_write_addr = 'd357;
        'd828 : mem_write_addr = 'd34;
        'd829 : mem_write_addr = 'd60;//
        'd830 : mem_write_addr = 'd117;
        'd831 : mem_write_addr = 'd269;
        'd832 : mem_write_addr = 'd164;
        'd833 : mem_write_addr = 'd186;
        'd834 : mem_write_addr = 'd207;
        'd835 : mem_write_addr = 'd339;
        'd836 : mem_write_addr = 'd35;
        'd837 : mem_write_addr = 'd61;
        'd838 : mem_write_addr = 'd118;
        'd839 : mem_write_addr = 'd270;// 
        'd840 : mem_write_addr = 'd165;
        'd841 : mem_write_addr = 'd187;
        'd842 : mem_write_addr = 'd320;
        'd843 : mem_write_addr = 'd36;
        'd844 : mem_write_addr = 'd62;
        'd845 : mem_write_addr = 'd119;
        'd846 : mem_write_addr = 'd271;
        'd847 : mem_write_addr = 'd166;
        'd848 : mem_write_addr = 'd188;
        'd849 : mem_write_addr = 'd37;// 
        'd850 : mem_write_addr = 'd63;
        'd851 : mem_write_addr = 'd120;
        'd852 : mem_write_addr = 'd144;
        'd853 : mem_write_addr = 'd167;
        'd854 : mem_write_addr = 'd38;
        'd855 : mem_write_addr = 'd80;
        'd856 : mem_write_addr = 'd121;
        'd857 : mem_write_addr = 'd145;
        'd858 : mem_write_addr = 'd39;
        'd859 : mem_write_addr = 'd81;// 
        'd860 : mem_write_addr = 'd122;
        'd861 : mem_write_addr = 'd40;
        'd862 : mem_write_addr = 'd82;
        'd863 : mem_write_addr = 'd41;
        default: mem_write_addr = 'd512;
    endcase
    
end
endmodule